package defines;

parameter SIZE_DATA = 8;

endpackage


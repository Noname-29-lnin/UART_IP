module Tx();

endmodule

module check_parity();

endmodule


module overrun();

endmodule

